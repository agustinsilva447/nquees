library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity top_nqueens is
generic(
        F : integer; -- depth of the fifo
        M : integer; -- size of the board MxM
        Q : integer; -- columns in pre-solution
        N : integer  -- N-1 bits required to count upto size of the board;
    );  
port(
    clk     : in  std_logic;
    p_nRst  : in  std_logic; 
    p_empt  : in  std_logic; 
    p_din   : in  std_logic_vector(31 downto 0);
    counter : out std_logic_vector(63 downto 0);
    done    : out std_logic;
    p_fread : out std_logic
    );
end entity;

architecture rtl of top_nqueens is 

    type array_out is array (M-1 downto 0) of std_logic_vector(N-1 downto 0); 
    signal asout_array: array_out; 

    constant K_19: integer := 19; 
    signal a_in_19: std_logic_vector((N*K_19-1) downto 0); 
    signal a_out_19: std_logic_vector((N*(K_19+1)-1) downto 0); 
    signal ack_in_19, next_in_19, ack_out_19, next_out_19: std_logic; 
    signal output_state_19: std_logic_vector(2 downto 0); 
    signal wen19, ren19, aful19, emp19: std_logic; 
    signal din19, dou19: std_logic_vector((N*K_19-1) downto 0); 

    constant K_18: integer := 18; 
    signal a_in_18: std_logic_vector((N*K_18-1) downto 0); 
    signal a_out_18: std_logic_vector((N*(K_18+1)-1) downto 0); 
    signal ack_in_18, next_in_18, ack_out_18, next_out_18: std_logic; 
    signal output_state_18: std_logic_vector(2 downto 0); 
    signal wen18, ren18, aful18, emp18: std_logic; 
    signal din18, dou18: std_logic_vector((N*K_18-1) downto 0); 

    constant K_17: integer := 17; 
    signal a_in_17: std_logic_vector((N*K_17-1) downto 0); 
    signal a_out_17: std_logic_vector((N*(K_17+1)-1) downto 0); 
    signal ack_in_17, next_in_17, ack_out_17, next_out_17: std_logic; 
    signal output_state_17: std_logic_vector(2 downto 0); 
    signal wen17, ren17, aful17, emp17: std_logic; 
    signal din17, dou17: std_logic_vector((N*K_17-1) downto 0); 

    constant K_16: integer := 16; 
    signal a_in_16: std_logic_vector((N*K_16-1) downto 0); 
    signal a_out_16: std_logic_vector((N*(K_16+1)-1) downto 0); 
    signal ack_in_16, next_in_16, ack_out_16, next_out_16: std_logic; 
    signal output_state_16: std_logic_vector(2 downto 0); 
    signal wen16, ren16, aful16, emp16: std_logic; 
    signal din16, dou16: std_logic_vector((N*K_16-1) downto 0); 

    constant K_15: integer := 15; 
    signal a_in_15: std_logic_vector((N*K_15-1) downto 0); 
    signal a_out_15: std_logic_vector((N*(K_15+1)-1) downto 0); 
    signal ack_in_15, next_in_15, ack_out_15, next_out_15: std_logic; 
    signal output_state_15: std_logic_vector(2 downto 0); 
    signal wen15, ren15, aful15, emp15: std_logic; 
    signal din15, dou15: std_logic_vector((N*K_15-1) downto 0); 

    constant K_14: integer := 14; 
    signal a_in_14: std_logic_vector((N*K_14-1) downto 0); 
    signal a_out_14: std_logic_vector((N*(K_14+1)-1) downto 0); 
    signal ack_in_14, next_in_14, ack_out_14, next_out_14: std_logic; 
    signal output_state_14: std_logic_vector(2 downto 0); 
    signal wen14, ren14, aful14, emp14: std_logic; 
    signal din14, dou14: std_logic_vector((N*K_14-1) downto 0); 

    constant K_13: integer := 13; 
    signal a_in_13: std_logic_vector((N*K_13-1) downto 0); 
    signal a_out_13: std_logic_vector((N*(K_13+1)-1) downto 0); 
    signal ack_in_13, next_in_13, ack_out_13, next_out_13: std_logic; 
    signal output_state_13: std_logic_vector(2 downto 0); 
    signal wen13, ren13, aful13, emp13: std_logic; 
    signal din13, dou13: std_logic_vector((N*K_13-1) downto 0); 

    constant K_12: integer := 12; 
    signal a_in_12: std_logic_vector((N*K_12-1) downto 0); 
    signal a_out_12: std_logic_vector((N*(K_12+1)-1) downto 0); 
    signal ack_in_12, next_in_12, ack_out_12, next_out_12: std_logic; 
    signal output_state_12: std_logic_vector(2 downto 0); 
    signal wen12, ren12, aful12, emp12: std_logic; 
    signal din12, dou12: std_logic_vector((N*K_12-1) downto 0); 

    constant K_11: integer := 11; 
    signal a_in_11: std_logic_vector((N*K_11-1) downto 0); 
    signal a_out_11: std_logic_vector((N*(K_11+1)-1) downto 0); 
    signal ack_in_11, next_in_11, ack_out_11, next_out_11: std_logic; 
    signal output_state_11: std_logic_vector(2 downto 0); 
    signal wen11, ren11, aful11, emp11: std_logic; 
    signal din11, dou11: std_logic_vector((N*K_11-1) downto 0); 

    constant K_10: integer := 10; 
    signal a_in_10: std_logic_vector((N*K_10-1) downto 0); 
    signal a_out_10: std_logic_vector((N*(K_10+1)-1) downto 0); 
    signal ack_in_10, next_in_10, ack_out_10, next_out_10: std_logic; 
    signal output_state_10: std_logic_vector(2 downto 0); 
    signal wen10, ren10, aful10, emp10: std_logic; 
    signal din10, dou10: std_logic_vector((N*K_10-1) downto 0); 

    constant K_9: integer := 9; 
    signal a_in_9: std_logic_vector((N*K_9-1) downto 0); 
    signal a_out_9: std_logic_vector((N*(K_9+1)-1) downto 0); 
    signal ack_in_9, next_in_9, ack_out_9, next_out_9: std_logic; 
    signal output_state_9: std_logic_vector(2 downto 0); 
    signal wen9, ren9, aful9, emp9: std_logic; 
    signal din9, dou9: std_logic_vector((N*K_9-1) downto 0); 

    constant K_8: integer := 8; 
    signal a_in_8: std_logic_vector((N*K_8-1) downto 0); 
    signal a_out_8: std_logic_vector((N*(K_8+1)-1) downto 0); 
    signal ack_in_8, next_in_8, ack_out_8, next_out_8: std_logic; 
    signal output_state_8: std_logic_vector(2 downto 0); 
    signal wen8, ren8, aful8, emp8: std_logic; 
    signal din8, dou8: std_logic_vector((N*K_8-1) downto 0); 

    constant K_7: integer := 7; 
    signal a_in_7: std_logic_vector((N*K_7-1) downto 0); 
    signal a_out_7: std_logic_vector((N*(K_7+1)-1) downto 0); 
    signal ack_in_7, next_in_7, ack_out_7, next_out_7: std_logic; 
    signal output_state_7: std_logic_vector(2 downto 0); 
    signal wen7, ren7, aful7, emp7: std_logic; 
    signal din7, dou7: std_logic_vector((N*K_7-1) downto 0); 

    constant K_6: integer := 6; 
    signal a_in_6: std_logic_vector((N*K_6-1) downto 0); 
    signal a_out_6: std_logic_vector((N*(K_6+1)-1) downto 0); 
    signal ack_in_6, next_in_6, ack_out_6, next_out_6: std_logic; 
    signal output_state_6: std_logic_vector(2 downto 0); 
    signal wen6, ren6, aful6, emp6: std_logic; 
    signal din6, dou6: std_logic_vector((N*K_6-1) downto 0); 

    constant K_5: integer := 5; 
    signal a_in_5: std_logic_vector((N*K_5-1) downto 0); 
    signal a_out_5: std_logic_vector((N*(K_5+1)-1) downto 0); 
    signal ack_in_5, next_in_5, ack_out_5, next_out_5: std_logic; 
    signal output_state_5: std_logic_vector(2 downto 0); 
    signal wen5, ren5, aful5, emp5: std_logic; 
    signal din5, dou5: std_logic_vector((N*K_5-1) downto 0); 

    constant K_4: integer := 4; 
    signal a_in_4: std_logic_vector((N*K_4-1) downto 0); 
    signal a_out_4: std_logic_vector((N*(K_4+1)-1) downto 0); 
    signal ack_in_4, next_in_4, ack_out_4, next_out_4: std_logic; 
    signal output_state_4: std_logic_vector(2 downto 0); 
    signal wen4, ren4, aful4, emp4: std_logic; 
    signal din4, dou4: std_logic_vector((N*K_4-1) downto 0); 

    constant K_3: integer := 3; 
    signal a_in_3: std_logic_vector((N*K_3-1) downto 0); 
    signal a_out_3: std_logic_vector((N*(K_3+1)-1) downto 0); 
    signal ack_in_3, next_in_3, ack_out_3, next_out_3: std_logic; 
    signal output_state_3: std_logic_vector(2 downto 0); 
    signal wen3, ren3, aful3, emp3: std_logic; 
    signal din3, dou3: std_logic_vector((N*K_3-1) downto 0); 

    constant K_2: integer := 2; 
    signal a_in_2: std_logic_vector((N*K_2-1) downto 0); 
    signal a_out_2: std_logic_vector((N*(K_2+1)-1) downto 0); 
    signal ack_in_2, next_in_2, ack_out_2, next_out_2: std_logic; 
    signal output_state_2: std_logic_vector(2 downto 0); 
    signal wen2, ren2, aful2, emp2: std_logic; 
    signal din2, dou2: std_logic_vector((N*K_2-1) downto 0); 

    signal s_nonzero: std_logic; 
    signal array_zeros: std_logic_vector(M-1 downto 0); 
    signal last_solu: std_logic_vector((N*(K_19+1)-1) downto 0); 
    signal last_candi: unsigned(N-1 downto 0); 
    signal last_digit: unsigned(N-1 downto 0); 
    signal counter_s: unsigned(63 downto 0); 
    signal nRst, done_s: std_logic; 
    signal fread, fempt: std_logic; 
    constant impar_vector: std_logic_vector(0 downto 0) := std_logic_vector(to_unsigned(M mod 2, 1)); 
    constant impar: std_logic := impar_vector(0);

      function f_BITWISE_AND ( 
        var_asout_array_1 : in std_logic_vector) 
        return std_logic is 
        variable v_AND: std_logic := '1'; 
      begin 
        for i in 0 to N-1 loop 
            v_AND := v_AND and (not var_asout_array_1(i)); 
        end loop; 
        return v_AND; 
      end function f_BITWISE_AND; 

      function f_BITWISE_OR ( 
        var_asout_array_2    : in std_logic_vector) 
        return std_logic is 
        variable v_OR : std_logic := '0'; 
      begin 
        for i in 0 to M-1 loop 
            v_OR := v_OR or var_asout_array_2(i); 
        end loop; 
        return v_OR; 
      end function f_BITWISE_OR; 

begin 

    fsm_19: entity work.fsm 
    generic map (K => 19, M => M, N =>N) 
    port map (clk=>clk, nRst=>nRst, a_in=>a_in_19, ack_in=>ack_in_19, next_in=>next_in_19, a_out=>a_out_19, ack_out=>ack_out_19, next_out=>next_out_19, output_state=>output_state_19); 

    fsm_18: entity work.fsm 
    generic map (K => 18, M => M, N =>N) 
    port map (clk=>clk, nRst=>nRst, a_in=>a_in_18, ack_in=>ack_in_18, next_in=>next_in_18, a_out=>a_out_18, ack_out=>ack_out_18, next_out=>next_out_18, output_state=>output_state_18); 

    fsm_17: entity work.fsm 
    generic map (K => 17, M => M, N =>N) 
    port map (clk=>clk, nRst=>nRst, a_in=>a_in_17, ack_in=>ack_in_17, next_in=>next_in_17, a_out=>a_out_17, ack_out=>ack_out_17, next_out=>next_out_17, output_state=>output_state_17); 

    fsm_16: entity work.fsm 
    generic map (K => 16, M => M, N =>N) 
    port map (clk=>clk, nRst=>nRst, a_in=>a_in_16, ack_in=>ack_in_16, next_in=>next_in_16, a_out=>a_out_16, ack_out=>ack_out_16, next_out=>next_out_16, output_state=>output_state_16); 

    fsm_15: entity work.fsm 
    generic map (K => 15, M => M, N =>N) 
    port map (clk=>clk, nRst=>nRst, a_in=>a_in_15, ack_in=>ack_in_15, next_in=>next_in_15, a_out=>a_out_15, ack_out=>ack_out_15, next_out=>next_out_15, output_state=>output_state_15); 

    fsm_14: entity work.fsm 
    generic map (K => 14, M => M, N =>N) 
    port map (clk=>clk, nRst=>nRst, a_in=>a_in_14, ack_in=>ack_in_14, next_in=>next_in_14, a_out=>a_out_14, ack_out=>ack_out_14, next_out=>next_out_14, output_state=>output_state_14); 

    fsm_13: entity work.fsm 
    generic map (K => 13, M => M, N =>N) 
    port map (clk=>clk, nRst=>nRst, a_in=>a_in_13, ack_in=>ack_in_13, next_in=>next_in_13, a_out=>a_out_13, ack_out=>ack_out_13, next_out=>next_out_13, output_state=>output_state_13); 

    fsm_12: entity work.fsm 
    generic map (K => 12, M => M, N =>N) 
    port map (clk=>clk, nRst=>nRst, a_in=>a_in_12, ack_in=>ack_in_12, next_in=>next_in_12, a_out=>a_out_12, ack_out=>ack_out_12, next_out=>next_out_12, output_state=>output_state_12); 

    fsm_11: entity work.fsm 
    generic map (K => 11, M => M, N =>N) 
    port map (clk=>clk, nRst=>nRst, a_in=>a_in_11, ack_in=>ack_in_11, next_in=>next_in_11, a_out=>a_out_11, ack_out=>ack_out_11, next_out=>next_out_11, output_state=>output_state_11); 

    fsm_10: entity work.fsm 
    generic map (K => 10, M => M, N =>N) 
    port map (clk=>clk, nRst=>nRst, a_in=>a_in_10, ack_in=>ack_in_10, next_in=>next_in_10, a_out=>a_out_10, ack_out=>ack_out_10, next_out=>next_out_10, output_state=>output_state_10); 

    fsm_9: entity work.fsm 
    generic map (K => 9, M => M, N =>N) 
    port map (clk=>clk, nRst=>nRst, a_in=>a_in_9, ack_in=>ack_in_9, next_in=>next_in_9, a_out=>a_out_9, ack_out=>ack_out_9, next_out=>next_out_9, output_state=>output_state_9); 

    fsm_8: entity work.fsm 
    generic map (K => 8, M => M, N =>N) 
    port map (clk=>clk, nRst=>nRst, a_in=>a_in_8, ack_in=>ack_in_8, next_in=>next_in_8, a_out=>a_out_8, ack_out=>ack_out_8, next_out=>next_out_8, output_state=>output_state_8); 

    fsm_7: entity work.fsm 
    generic map (K => 7, M => M, N =>N) 
    port map (clk=>clk, nRst=>nRst, a_in=>a_in_7, ack_in=>ack_in_7, next_in=>next_in_7, a_out=>a_out_7, ack_out=>ack_out_7, next_out=>next_out_7, output_state=>output_state_7); 

    fsm_6: entity work.fsm 
    generic map (K => 6, M => M, N =>N) 
    port map (clk=>clk, nRst=>nRst, a_in=>a_in_6, ack_in=>ack_in_6, next_in=>next_in_6, a_out=>a_out_6, ack_out=>ack_out_6, next_out=>next_out_6, output_state=>output_state_6); 

    fsm_5: entity work.fsm 
    generic map (K => 5, M => M, N =>N) 
    port map (clk=>clk, nRst=>nRst, a_in=>a_in_5, ack_in=>ack_in_5, next_in=>next_in_5, a_out=>a_out_5, ack_out=>ack_out_5, next_out=>next_out_5, output_state=>output_state_5); 

    fsm_4: entity work.fsm 
    generic map (K => 4, M => M, N =>N) 
    port map (clk=>clk, nRst=>nRst, a_in=>a_in_4, ack_in=>ack_in_4, next_in=>next_in_4, a_out=>a_out_4, ack_out=>ack_out_4, next_out=>next_out_4, output_state=>output_state_4); 

    fsm_3: entity work.fsm 
    generic map (K => 3, M => M, N =>N) 
    port map (clk=>clk, nRst=>nRst, a_in=>a_in_3, ack_in=>ack_in_3, next_in=>next_in_3, a_out=>a_out_3, ack_out=>ack_out_3, next_out=>next_out_3, output_state=>output_state_3); 

    fsm_2: entity work.fsm 
    generic map (K => 2, M => M, N =>N) 
    port map (clk=>clk, nRst=>nRst, a_in=>a_in_2, ack_in=>ack_in_2, next_in=>next_in_2, a_out=>a_out_2, ack_out=>ack_out_2, next_out=>next_out_2, output_state=>output_state_2); 

    fifo_19: entity work.fifo 
    generic map(DWIDTH => N*K_19, DEPTH => F, AFULLOFFSET => 1, AEMPTYOFFSET => 1, ASYNC => False) 
    port map(wclk_i=>clk, rclk_i=>clk, wrst_i=>nRst, rrst_i=>nRst, data_i => din19, wen_i => wen19, ren_i => ren19, data_o => dou19, afull_o => aful19, empty_o => emp19); 

    fifo_18: entity work.fifo 
    generic map(DWIDTH => N*K_18, DEPTH => F, AFULLOFFSET => 1, AEMPTYOFFSET => 1, ASYNC => False) 
    port map(wclk_i=>clk, rclk_i=>clk, wrst_i=>nRst, rrst_i=>nRst, data_i => din18, wen_i => wen18, ren_i => ren18, data_o => dou18, afull_o => aful18, empty_o => emp18); 

    fifo_17: entity work.fifo 
    generic map(DWIDTH => N*K_17, DEPTH => F, AFULLOFFSET => 1, AEMPTYOFFSET => 1, ASYNC => False) 
    port map(wclk_i=>clk, rclk_i=>clk, wrst_i=>nRst, rrst_i=>nRst, data_i => din17, wen_i => wen17, ren_i => ren17, data_o => dou17, afull_o => aful17, empty_o => emp17); 

    fifo_16: entity work.fifo 
    generic map(DWIDTH => N*K_16, DEPTH => F, AFULLOFFSET => 1, AEMPTYOFFSET => 1, ASYNC => False) 
    port map(wclk_i=>clk, rclk_i=>clk, wrst_i=>nRst, rrst_i=>nRst, data_i => din16, wen_i => wen16, ren_i => ren16, data_o => dou16, afull_o => aful16, empty_o => emp16); 

    fifo_15: entity work.fifo 
    generic map(DWIDTH => N*K_15, DEPTH => F, AFULLOFFSET => 1, AEMPTYOFFSET => 1, ASYNC => False) 
    port map(wclk_i=>clk, rclk_i=>clk, wrst_i=>nRst, rrst_i=>nRst, data_i => din15, wen_i => wen15, ren_i => ren15, data_o => dou15, afull_o => aful15, empty_o => emp15); 

    fifo_14: entity work.fifo 
    generic map(DWIDTH => N*K_14, DEPTH => F, AFULLOFFSET => 1, AEMPTYOFFSET => 1, ASYNC => False) 
    port map(wclk_i=>clk, rclk_i=>clk, wrst_i=>nRst, rrst_i=>nRst, data_i => din14, wen_i => wen14, ren_i => ren14, data_o => dou14, afull_o => aful14, empty_o => emp14); 

    fifo_13: entity work.fifo 
    generic map(DWIDTH => N*K_13, DEPTH => F, AFULLOFFSET => 1, AEMPTYOFFSET => 1, ASYNC => False) 
    port map(wclk_i=>clk, rclk_i=>clk, wrst_i=>nRst, rrst_i=>nRst, data_i => din13, wen_i => wen13, ren_i => ren13, data_o => dou13, afull_o => aful13, empty_o => emp13); 

    fifo_12: entity work.fifo 
    generic map(DWIDTH => N*K_12, DEPTH => F, AFULLOFFSET => 1, AEMPTYOFFSET => 1, ASYNC => False) 
    port map(wclk_i=>clk, rclk_i=>clk, wrst_i=>nRst, rrst_i=>nRst, data_i => din12, wen_i => wen12, ren_i => ren12, data_o => dou12, afull_o => aful12, empty_o => emp12); 

    fifo_11: entity work.fifo 
    generic map(DWIDTH => N*K_11, DEPTH => F, AFULLOFFSET => 1, AEMPTYOFFSET => 1, ASYNC => False) 
    port map(wclk_i=>clk, rclk_i=>clk, wrst_i=>nRst, rrst_i=>nRst, data_i => din11, wen_i => wen11, ren_i => ren11, data_o => dou11, afull_o => aful11, empty_o => emp11); 

    fifo_10: entity work.fifo 
    generic map(DWIDTH => N*K_10, DEPTH => F, AFULLOFFSET => 1, AEMPTYOFFSET => 1, ASYNC => False) 
    port map(wclk_i=>clk, rclk_i=>clk, wrst_i=>nRst, rrst_i=>nRst, data_i => din10, wen_i => wen10, ren_i => ren10, data_o => dou10, afull_o => aful10, empty_o => emp10); 

    fifo_9: entity work.fifo 
    generic map(DWIDTH => N*K_9, DEPTH => F, AFULLOFFSET => 1, AEMPTYOFFSET => 1, ASYNC => False) 
    port map(wclk_i=>clk, rclk_i=>clk, wrst_i=>nRst, rrst_i=>nRst, data_i => din9, wen_i => wen9, ren_i => ren9, data_o => dou9, afull_o => aful9, empty_o => emp9); 

    fifo_8: entity work.fifo 
    generic map(DWIDTH => N*K_8, DEPTH => F, AFULLOFFSET => 1, AEMPTYOFFSET => 1, ASYNC => False) 
    port map(wclk_i=>clk, rclk_i=>clk, wrst_i=>nRst, rrst_i=>nRst, data_i => din8, wen_i => wen8, ren_i => ren8, data_o => dou8, afull_o => aful8, empty_o => emp8); 

    fifo_7: entity work.fifo 
    generic map(DWIDTH => N*K_7, DEPTH => F, AFULLOFFSET => 1, AEMPTYOFFSET => 1, ASYNC => False) 
    port map(wclk_i=>clk, rclk_i=>clk, wrst_i=>nRst, rrst_i=>nRst, data_i => din7, wen_i => wen7, ren_i => ren7, data_o => dou7, afull_o => aful7, empty_o => emp7); 

    fifo_6: entity work.fifo 
    generic map(DWIDTH => N*K_6, DEPTH => F, AFULLOFFSET => 1, AEMPTYOFFSET => 1, ASYNC => False) 
    port map(wclk_i=>clk, rclk_i=>clk, wrst_i=>nRst, rrst_i=>nRst, data_i => din6, wen_i => wen6, ren_i => ren6, data_o => dou6, afull_o => aful6, empty_o => emp6); 

    fifo_5: entity work.fifo 
    generic map(DWIDTH => N*K_5, DEPTH => F, AFULLOFFSET => 1, AEMPTYOFFSET => 1, ASYNC => False) 
    port map(wclk_i=>clk, rclk_i=>clk, wrst_i=>nRst, rrst_i=>nRst, data_i => din5, wen_i => wen5, ren_i => ren5, data_o => dou5, afull_o => aful5, empty_o => emp5); 

    fifo_4: entity work.fifo 
    generic map(DWIDTH => N*K_4, DEPTH => F, AFULLOFFSET => 1, AEMPTYOFFSET => 1, ASYNC => False) 
    port map(wclk_i=>clk, rclk_i=>clk, wrst_i=>nRst, rrst_i=>nRst, data_i => din4, wen_i => wen4, ren_i => ren4, data_o => dou4, afull_o => aful4, empty_o => emp4); 

    fifo_3: entity work.fifo 
    generic map(DWIDTH => N*K_3, DEPTH => F, AFULLOFFSET => 1, AEMPTYOFFSET => 1, ASYNC => False) 
    port map(wclk_i=>clk, rclk_i=>clk, wrst_i=>nRst, rrst_i=>nRst, data_i => din3, wen_i => wen3, ren_i => ren3, data_o => dou3, afull_o => aful3, empty_o => emp3); 

    fifo_2: entity work.fifo 
    generic map(DWIDTH => N*K_2, DEPTH => F, AFULLOFFSET => 1, AEMPTYOFFSET => 1, ASYNC => False) 
    port map(wclk_i=>clk, rclk_i=>clk, wrst_i=>nRst, rrst_i=>nRst, data_i => din2, wen_i => wen2, ren_i => ren2, data_o => dou2, afull_o => aful2, empty_o => emp2); 

    ack_in_19 <= emp19; 
    a_in_19 <= dou19; 
    ren19 <= next_out_19; 
    wen19 <= not ack_out_18; 
    din19 <= a_out_18; 
    next_in_18 <= not aful19; 

    ack_in_18 <= emp18; 
    a_in_18 <= dou18; 
    ren18 <= next_out_18; 
    wen18 <= not ack_out_17; 
    din18 <= a_out_17; 
    next_in_17 <= not aful18; 

    ack_in_17 <= emp17; 
    a_in_17 <= dou17; 
    ren17 <= next_out_17; 
    wen17 <= not ack_out_16; 
    din17 <= a_out_16; 
    next_in_16 <= not aful17; 

    ack_in_16 <= emp16; 
    a_in_16 <= dou16; 
    ren16 <= next_out_16; 
    wen16 <= not ack_out_15; 
    din16 <= a_out_15; 
    next_in_15 <= not aful16; 

    ack_in_15 <= emp15; 
    a_in_15 <= dou15; 
    ren15 <= next_out_15; 
    wen15 <= not ack_out_14; 
    din15 <= a_out_14; 
    next_in_14 <= not aful15; 

    ack_in_14 <= emp14; 
    a_in_14 <= dou14; 
    ren14 <= next_out_14; 
    wen14 <= not ack_out_13; 
    din14 <= a_out_13; 
    next_in_13 <= not aful14; 

    ack_in_13 <= emp13; 
    a_in_13 <= dou13; 
    ren13 <= next_out_13; 
    wen13 <= not ack_out_12; 
    din13 <= a_out_12; 
    next_in_12 <= not aful13; 

    ack_in_12 <= emp12; 
    a_in_12 <= dou12; 
    ren12 <= next_out_12; 
    wen12 <= not ack_out_11; 
    din12 <= a_out_11; 
    next_in_11 <= not aful12; 

    ack_in_11 <= emp11; 
    a_in_11 <= dou11; 
    ren11 <= next_out_11; 
    wen11 <= not ack_out_10; 
    din11 <= a_out_10; 
    next_in_10 <= not aful11; 

    ack_in_10 <= emp10; 
    a_in_10 <= dou10; 
    ren10 <= next_out_10; 
    wen10 <= not ack_out_9; 
    din10 <= a_out_9; 
    next_in_9 <= not aful10; 

    ack_in_9 <= emp9; 
    a_in_9 <= dou9; 
    ren9 <= next_out_9; 
    wen9 <= not ack_out_8; 
    din9 <= a_out_8; 
    next_in_8 <= not aful9; 

    ack_in_8 <= emp8; 
    a_in_8 <= dou8; 
    ren8 <= next_out_8; 
    wen8 <= not ack_out_7; 
    din8 <= a_out_7; 
    next_in_7 <= not aful8; 

    ack_in_7 <= emp7; 
    a_in_7 <= dou7; 
    ren7 <= next_out_7; 
    wen7 <= not ack_out_6; 
    din7 <= a_out_6; 
    next_in_6 <= not aful7; 

    ack_in_6 <= emp6; 
    a_in_6 <= dou6; 
    ren6 <= next_out_6; 
    wen6 <= not ack_out_5; 
    din6 <= a_out_5; 
    next_in_5 <= not aful6; 

    ack_in_5 <= emp5; 
    a_in_5 <= dou5; 
    ren5 <= next_out_5; 
    wen5 <= not ack_out_4; 
    din5 <= a_out_4; 
    next_in_4 <= not aful5; 

    ack_in_4 <= emp4; 
    a_in_4 <= dou4; 
    ren4 <= next_out_4; 
    wen4 <= not ack_out_3; 
    din4 <= a_out_3; 
    next_in_3 <= not aful4; 

    ack_in_3 <= emp3; 
    a_in_3 <= dou3; 
    ren3 <= next_out_3; 
    wen3 <= not ack_out_2; 
    din3 <= a_out_2; 
    next_in_2 <= not aful3; 

    ack_in_2 <= emp2; 
    a_in_2 <= dou2; 
    ren2 <= next_out_2; 
    done <= done_s; 
    nRst <= p_nRst; 
    counter <= std_logic_vector(counter_s); 
    last_digit <= unsigned(a_in_19((N*(M-1)-1) downto (N*(M-2)))); 
    last_candi <= (to_unsigned(M/2, N) + 1)  when impar = '1' else 
                  (to_unsigned(M/2, N))      when impar = '0'; 

    din2   <= p_din(N*Q-1 downto 0); 
    fempt   <= p_empt; 
    wen2    <= fread; 
    p_fread <= fread; 

    GENERATE_FOR_out: for i in 0 to M-1 generate 
        asout_array(i) <= a_out_19((N*(i+1)-1) downto N*i); 
    end generate;         
    GENERATE_FOR_zeros: for i in 0 to M-1 generate 
        array_zeros(i) <= f_BITWISE_AND(asout_array(i)); 
    end generate; 
    s_nonzero   <= f_BITWISE_OR(array_zeros); 
 
    counter_process: process(nRst, clk) 
    begin 
        if nRst = '1' then 
            next_in_19 <= '0'; 
            counter_s <= (others=>'0'); 
            last_solu <= (others=>'0'); 
        else 
            next_in_19 <= '1'; 
            if (clk'event and clk = '1') then 
                if (ack_out_19 = '0' and s_nonzero = '0' and last_solu /= a_out_19) then 
                    last_solu <= a_out_19; 
                    if (impar = '1' and last_digit = last_candi) then 
                        counter_s <= counter_s + 1; 
                    else 
                        counter_s <= counter_s + 2; 
                    end if; 
                end if; 
            end if; 
        end if; 
    end process; 

    reading_process: process(nRst, clk) 
    begin 
        if nRst = '1' then 
            done_s <= '0'; 
            fread <= '0'; 
        elsif (clk'event and clk = '1') then 
            done_s <= (emp2 and emp3 and emp4 and emp5 and emp6 and emp7 and emp8 and emp9 and emp10 and emp11 and emp12 and emp13 and emp14 and emp15 and emp16 and emp17 and emp18 and emp19); 
            if (fempt = '0' and aful2 = '0') then 
                fread <= '1'; 
            else 
                fread <= '0'; 
            end if; 
        end if; 
    end process; 

end architecture;